

module hw1test;
reg A; // inputs 
reg B;

wire nA; // intermediate wires
wire nB;
wire nAandnB;
wire AandB;
wire nAandB;
wire nAornB;
wire AorB;
wire nAorB;

// ~(AB)
and one(AandB, A, B);
not two(nAandB, AandB);

// (~A)+(~B)
not thee(nA, A);
not four(nB, B);
or five(nAornB, nA, nB);

// ~(A+B)
or six(AorB, A, B);
not seven(nAorB, AorB);

// (~A)(~B)
not eight(nA, A);
not nine(nB, B);
and ten(nAandnB, nA, nB);



initial begin
$display("A B | ~A ~B | ~(AB) ~A+~B | ~(A+B) ~A~B");
A=0;B=0; #1
$display("%b %b |  %b  %b |    %b    %b   |    %b    %b", A,B, nA, nB, nAandB, nAornB, nAorB, nAandnB);
A=0; B=1; #1
$display("%b %b |  %b  %b |    %b    %b   |    %b    %b", A,B, nA, nB, nAandB, nAornB, nAorB, nAandnB);
A=1; B=0; #1
$display("%b %b |  %b  %b |    %b    %b   |    %b    %b", A,B, nA, nB, nAandB, nAornB, nAorB, nAandnB);
A=1; B=1; #1
$display("%b %b |  %b  %b |    %b    %b   |    %b    %b", A,B, nA, nB, nAandB, nAornB, nAorB, nAandnB);

end

endmodule;
